module NAND
(
  input logic a, b,
  output logic y
);
  assign y = ~(a & b);
endmodule
